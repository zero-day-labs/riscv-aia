`define MSI_MODE
// `define DIRECT_MODE